module 7SegmentDecoder #(parameter WIDTH = 4) (
    input [WIDTH-1:0] b,
    output [6:0] c,
[6:0] c = 0;
if(b == 0)(//0
    [6:0] c = [1 0 0 0 0 0 0];
)
if(b==[0 0 0 1])(//1
    [6:0] c = [1 1 1 1 0 0 1];
)
if(b==[0 0 1 0])(//2
    [6:0] c = [0 1 0 0 1 0 0];
)
if(b==[0 0 1 1])(//3
    [6:0] c = [0 1 1 0 0 0 0];
)
if(b==[0 1 0 0])(//4
    [6:0] c = [0 0 1 1 0 0 1];
)
if(b==[0 1 0 1])(//5
    [6:0] c = [0 0 1 0 0 1 0];
)
if(b==[0 1 1 0])(//6
    [6:0] c = [0 0 0 0 0 1 0];
)
if(b==[0 1 1 1])(//7
    [6:0] c = [1 1 1 1 0 0 0];
)
if(b==[1 0 0 0])(//8
    [6:0] c = [0 0 0 0 0 0 0];
)
if(b==[1 0 0 1])(//9
    [6:0] c = [0 0 1 0 0 0 0];
)
if(b==[1 0 1 0])(//A
    [6:0] c = [0 0 0 1 0 0 0];
)
if(b==[1 0 1 1])(//b
    [6:0] c = [0 0 0 0 0 1 1];
)
if(b==[1 1 0 0])(//C
    [6:0] c = [1 0 0 0 1 1 0];
)
if(b==[1 1 0 1])(//d
    [6:0] c = [0 1 0 0 0 0 1];
)
if(b==[1 1 1 0])(//E
    [6:0] c = [0 0 0 0 1 1 0];
)
if(b==[1 1 1 1])(//F
    [6:0] c = [0 0 0 1 1 1 0];
)
);
endmodule;